
module fpga_top_level(
	input reset,
	input clock,
	input [7:0]  writedata,
	input write,
	input chipselect,
	input [3:0]  address
);

	//vga_display vga_disp();
	//sdram_controller sdram_ctrl();

endmodule
