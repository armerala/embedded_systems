
module sdram_controller(
	input [14:0] mem_a,
	input [2:0] mem_ba,
	input mem_cas_n,
	input mem_ck,
	input mem_ck_n,
	input mem_cke,
	input mem_cs_n,
	input [3:0] mem_dm,
	input [31:0] mem_dq,
	input [3:0] mem_dqs,
	input [3:0] mem_dqs_n,
	input mem_odt,
	input mem_ras_n,
	input mem_reset_n,
	input mem_we_n,
	output oct_rzqin
);


endmodule
